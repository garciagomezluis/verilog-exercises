module greater_than_v2(input [1:0] A, input [1:0] B, output F);
    assign F = A > B;
endmodule
